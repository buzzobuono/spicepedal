.title Fender Bassman Tone Stack

R1 1 4 56k
C1 1 2 250e-12
C2 4 5 0.02e-6
Ptreble 2 5 3 250k param=treble Taper=LIN
W 5 6
Pbass 5 7 6 1M param=bass Taper=LIN
C3 4 8 0.02e-6
Pmid 7 0 8 25k param=mid Taper=LIN

.input 1 Z=50k
.output 3
.param bass 0.5
.param mid 0.5
.param treble 0.5
.ctrl 0 bass 0.0 1.0 0.1
.ctrl 1 mid 0.0 1.0 0.1
.ctrl 2 treble 0.0 1.0 0.1
.probe V(1) V(3)