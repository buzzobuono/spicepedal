.title Non-Inverting Summing Amplifier

VCC 10 0 DC 15
VEE 11 0 DC -15

* Due ingressi
V1 1 0 SIN(0 0.5 440)
V2 4 0 SIN(0 0.5 660)

* Somma passiva in ingresso
R1 1 2 10k
R2 4 2 10k

* Amplificatore non invertente
Rin 3 0 10k
Rf 3 2 20k

* OpAmp: output = node 3
XOP 3 2 3 10 11 OPAMP

.control
tran 0.1ms 5ms
plot v(1) v(4) v(3)
.endc
.end
