* Tremolo

B_LFO 0 0 Rs=1 V="modulation:=(depth * sin(2 * 3.14 * speed * t))"
B_GAIN 2 0 V="V(1) * (1 + modulation)" Rs=1

.param speed 8
.param depth 0.8
.param modulation 0
.input 1
.output 2
.probe tremolo.csv V(1) V(2)