.title Woolly Mammoth

VCC 9 0 DC 9

* two stage amplifier

R3 9 1 51k
R4 9 2 20k
Q1 1 3 0 Q2N3904
*Q2 2 1 5 Q2N3904
Q2.1 2 1 15 QMOD ; MPSA13
Q2.2 2 15 5 QMOD
.model QMOD Q Is=360f Bf=337 Br=4
.model 2N3904 Q Bf=160.1 Br=5.944 Is=4.639e-15 Vt=0.02585

R2 3 4 100k
Ppinch 4 5 8 500k param=pinch taper=LIN
W1 8 5

C6 5 6 100u
R1 8 0 2.2k
Pwool 6 11 0 2k param=wool taper=LIN

C1 7 3 0.22u
C2 3 0 10n

* tone stack

C3 2 10 10n
C5 2 11 100u
R5 11 10 10k
R5b 11 10 15k

R6 11 12 5.1k
C4 12 0 7.4n
C4b 12 0 220n

Peq 12 10 13 10k param=eq taper=LIN
Pvol 13 0 14 10k param=volume taper=LIN




.input 7
.output 14
.warmup 60
.param pinch .8
.param wool .8
.param eq .8
.param volume .8
.ctrl 0 pinch 0 1
.ctrl 1 wool 0 1
.ctrl 2 eq 0 1
.ctrl 3 volume 0 1
*.probe V(14)