.title Full Wave Rectifier

VCC 10 0 DC 15
VEE 11 0 DC -15

* Percorso diretto per semionda positiva
D1 1 2 1N4148
*D1 1 2 Schottky
Rload 2 0 50k

* Percorso invertente per semionda negativa
Rin 1 3 10k
Rf 3 4 10k
OP 4 0 3 10 11 TL072 Rout=75 Imax=0.020 Gain=10000 Sr=13

D2 4 2 1N4148
*D2 4 2 SchottkyInLine Is=1e-6 N=1.21 Vt=0.02585 Cj0=1e-12 Vj=0.3 Mj=0.02

* Carico finale
Rload2 2 0 50k

.model Schottky D Is=1e-7 N=1.1 Vt=0.02585 Cj0=1e-11 Vj=0.3 Mj=0.02
.include circuits/models/diodes.lib
.input 1
.output 2
.probe full-wave-rectifier.csv V(1) V(2)
