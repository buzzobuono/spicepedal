.title SHO booster
.param volume = 0.5


V1 0 1 -9
D1 3 1 D1N4148
D1 0 3 D1N4148
C1 in 3 0.1u
R3 1 2 5.1k
xQ1 2 3 4 BS170
R2 2 3 10m
R1 3 0 10m
C2 2 out 10u
XPOTVOLUME 4 0 0 POT PARAMS: VALUE=5K SET={volume}
R5 out 0 100k





.include "../../mylib.lib"

.model filesrc filesource (file="../../input/input.data" amploffset=[0] amplscale=[1]
+                          timeoffset=0 timescale=1
+                          timerelative=false amplstep=false)

.model D1N4148 D(IS=0.1P RS=16 CJO=2P TT=12N BV=100 IBV=0.1P)

.SUBCKT BS170 1 2 3
* 1=drain  2=gate  3=source
Cgs  2 3 12.3E-12
Cgd1 2 4 27.4E-12
Cgd2 1 4 6E-12
M1 1 2 3 3 MOST1
M2 4 2 1 3 MOST2
D1 3 1 Dbody
.MODEL MOST1 NMOS(Level=3 Kp=20.78u W=9.7m L=2u Rs=20m Vto=2 Rd=1.186)
.MODEL MOST2 NMOS(VTO=-4.73 Kp=20.78u W=9.7m L=2u Rs=20m)
.MODEL Dbody D(Is=125f N=1.023 Rs=1.281 Ikf=18.01 Cjo=46.3p M=.3423
+            Vj=.4519 Bv=60 Ibv=10u Tt=161.6n)
.ENDS

.INPUT
.OUTPUT