.title Convertitore Sinusoidale a Onda Quadra - Output 0.2V con partitore

VCC 10 0 DC 5
VEE 11 0 DC -5

* Amplificatore non invertente con guadagno elevato per saturazione
* Guadagno = 1 + R2/R1 = 1 + 90k/1k = 91
O1 3 1 2 10 11 TL072 Rout=75 Imax=0.020 Gain=10000 Sr=13

R1 2 0 1k
R2 3 2 90k

* Partitore resistivo per ridurre output da ±5V a ±0.2V
* Fattore di divisione = 0.2/5 = 0.04 = 1/25
R3 3 4 24k
R4 4 0 1k

.input 1
.output 4
* OpAmps
.model TL072 O Rout=75 Imax=0.020 Gain=10000 Sr=13
* 
.probe opamp-98-square-wave.csv V(input) V(1) V(4)
