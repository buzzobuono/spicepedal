.title Bazz Fuss

V1 1 0 DC 9
R1 1 2 100k
D1 2 3 D1N914
C2 2 4 0.1u
Q1 2 3 0 2N5088
*Q1 2 3 0 BC549BP
*Q1 2 3 0 NPN Bf=200 Br=1 Is=1e-14 Vt=0.026
C1 5 3 4.7u
R2 4 0 100M

Pvol0 4 0 7 100k param=volume taper=LOG

.input 5
.output 7
.include circuits/models/diodes.lib
.include circuits/models/transistors.lib
.probe V(5) V(7)
.ic C1 0.60683
.ic C2 0.50573
.warmup 2
.param volume 0.5
.ctrl 0 volume 0.0 1.0